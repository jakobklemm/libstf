`timescale 1ns / 1ps

`include "libstf_macros.svh"

/**
 * Converts an ndata_i stream to a different width.
 *
 * 8->16 & 16->8 supported
 */
module NDataWidthConverter #(
    parameter type data_t,
    parameter IN_WIDTH,
    parameter OUT_WIDTH
) (
    input logic clk,
    input logic rst_n,

    ndata_i.s in, // #(data_t, IN_WIDTH)
    ndata_i.m out // #(data_t, OUT_WIDTH)
);

generate if (IN_WIDTH == OUT_WIDTH) begin

`DATA_ASSIGN(in, out)

end else if (IN_WIDTH == 8 && OUT_WIDTH == 16) begin
    // 8 -> 16 conversion 

    logic is_upper, n_is_upper;

    data_t[OUT_WIDTH - 1:0] data,  n_data;
    logic[OUT_WIDTH - 1:0]  keep,  n_keep;
    logic                   last,  n_last;
    logic                   valid, n_valid;

    assign in.ready = out.ready;

    always_ff @(posedge clk) begin
        if (rst_n == 1'b0) begin
            is_upper <= 1'b0;

            valid <= 1'b0;
        end else begin
            is_upper <= n_is_upper;

            data  <= n_data;
            keep  <= n_keep;
            last  <= n_last;
            valid <= n_valid;
        end
    end

    always_comb begin
        n_is_upper = is_upper;

        n_data  = data;
        n_keep  = keep;
        n_last  = last;
        n_valid = 1'b0;

        if (out.ready) begin
            if (in.valid) begin
                if (!in.last) begin
                    n_is_upper = ~is_upper;
                end else begin
                    n_is_upper = 1'b0;
                end
            end

            if (!is_upper) begin
                n_data[7:0]  = in.data;
                n_keep[15:8] = '0;
                n_keep[7:0]  = in.keep;
                if (in.last) begin
                    n_valid = in.valid;
                end
            end else begin
                n_data[15:8] = in.data;
                n_keep[15:8] = in.keep;
                n_valid      = in.valid;
            end

            n_last = in.last;
        end else begin
            n_valid = valid;
        end
    end

    assign out.data  = data;
    assign out.keep  = keep;
    assign out.last  = last;
    assign out.valid = valid;

end else if (IN_WIDTH == 16 && OUT_WIDTH == 8) begin
    // 16 -> 8 conversion
    logic has_upper, n_has_upper;
    data_t[OUT_WIDTH - 1:0] upper_data,  n_upper_data;
    logic[OUT_WIDTH - 1:0]  upper_keep,  n_upper_keep;
    logic                   upper_last,  n_upper_last;

    always_ff @(posedge clk) begin
        if (rst_n == 1'b0) begin
            has_upper <= 1'b0;
        end else begin
            has_upper <= n_has_upper;
            upper_data  <= n_upper_data;
            upper_keep  <= n_upper_keep;
            upper_last  <= n_upper_last;
        end
    end

    always_comb begin
        n_has_upper = has_upper;
        n_upper_data = upper_data;
        n_upper_keep = upper_keep;
        n_upper_last = upper_last;

        if (out.ready && has_upper) begin
            // Output stored upper
            n_has_upper = 1'b0;
        end else if (in.valid && !has_upper && out.ready) begin
            // input is valid => output lower half, store upper half for next cycle
            n_has_upper = 1'b1;
            n_upper_data = in.data[15:8];
            n_upper_keep = in.keep[15:8];
            n_upper_last = in.last;
        end 
    end

    assign in.ready = out.ready && !has_upper;

    assign out.data  = has_upper ? upper_data : in.data[7:0];
    assign out.keep  = has_upper ? upper_keep : in.keep[7:0];
    assign out.last  = has_upper & upper_last;

    assign out.valid = has_upper || in.valid;

end else begin
    initial $error("NDataWidthConverter: unsupported");
end endgenerate

endmodule
